module DECODER(
    input [5:0] ins_op,
    output reg_write,
    output reg_dst,
    output alu_src,
    output pc_src,
    output [1:0] alu_op,
    output mem_read,
    output mem_write,
    output mem_to_reg
);


endmodule
